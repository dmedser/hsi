module hsi_s_tx_ctrl (
	input clk,
	input clk_en,
	input n_rst,
	input sd_busy,
	input sr,
	output dat1,
	output dat2
);

endmodule