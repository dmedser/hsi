/********** МАРКЕРЫ **********/
`define MARKER_MASTER 8'hA5
`define MARKER_SLAVE  8'hB6 

/*********** ФЛАГИ ***********/
`define FLAG_BOARD_TIME_CODE 		 8'h01
`define FLAG_CONTROL_COMMAND_WORD 8'h02
`define FLAG_STATUS_REQUEST 		 8'h03
`define FLAG_DATA_PACKET_REQUEST  8'h04
`define FLAG_TIME_MARK  			 8'h05
