`define SYS_TIME_REG_ADDR 	8'h00
`define SDI_CTRL_REG_ADDR 	8'h08
`define CSI_CTRL_REG_ADDR 	8'h0A
`define CCW_BUF_ADDR  		8'h0C
